`ifndef HBM_MANYCORE_VH
`define HBM_MANYCORE_VH

  `define USE_IP_GEN

  `define FPGA_LESS_RST

`endif
