`ifndef BSG_BLADERUNNER_DEFINES_VH
`define BSG_BLADERUNNER_DEFINES_VH

`define FPGA_TARGET_ULTRASCALE_PLUS

`endif
