/*
* qcl_dff_reset.v
*
*/

module qcl_dff_reset #(
  parameter width_p = 1
  , parameter reset_val_p = 0
) (
  input                clk_i
  ,input                reset_i
  ,input  [width_p-1:0] data_i
  ,output [width_p-1:0] data_o
);


`ifdef FPGA_LESS_RST
  logic [width_p-1:0] data_r = width_p'(reset_val_p);
`else
  logic [width_p-1:0] data_r;
`endif

  assign data_o = data_r;

  always_ff @(posedge clk_i) begin
    if (reset_i)
      data_r <= width_p'(reset_val_p);
    else
      data_r <= data_i;
  end

endmodule
