`ifndef BSG_BLADERUNNER_DEFINES_VH
`define BSG_BLADERUNNER_DEFINES_VH

`define FPGA_TARGET_ULTRASCALE_PLUS

`define FPGA_TARGET_HBM

`define FPGA_LESS_RST

`define USE_IP_GEN

`endif
